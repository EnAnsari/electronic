** Profile: "SCHEMATIC1-Y"  [ C:\Users\WOLF2022\Desktop\UNI\3_semiterm\MadarElectric\Az\word\10\Pr01\r-SCHEMATIC1-Y.sim ] 

** Creating circuit file "r-SCHEMATIC1-Y.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 10u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\r-SCHEMATIC1.net" 


.END
