** Profile: "SCHEMATIC1-T"  [ C:\Users\WOLF2022\Desktop\UNI\3_semiterm\MadarElectric\Az\word\13\TEST\t-schematic1-t.sim ] 

** Creating circuit file "t-schematic1-t.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 1 100meg
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\t-SCHEMATIC1.net" 


.END
