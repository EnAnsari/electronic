** Profile: "SCHEMATIC1-RL2"  [ C:\Users\WOLF2022\Desktop\UNI\3_semiterm\MadarElectric\Az\word\7\RL\rl-schematic1-rl2.sim ] 

** Creating circuit file "rl-schematic1-rl2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rl-SCHEMATIC1.net" 


.END
