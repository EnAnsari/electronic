** Profile: "SCHEMATIC1-th"  [ C:\Users\WOLF2022\Desktop\UNI\3_semiterm\MadarElectric\Az\word\4\thevenin\thevenin-SCHEMATIC1-th.sim ] 

** Creating circuit file "thevenin-SCHEMATIC1-th.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\thevenin-SCHEMATIC1.net" 


.END
