** Profile: "SCHEMATIC1-Rec"  [ C:\Users\WOLF2022\Desktop\UNI\3_semiterm\MadarElectric\Az\word\10\Pr\rectifire-schematic1-rec.sim ] 

** Creating circuit file "rectifire-schematic1-rec.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1s 0 1000u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rectifire-SCHEMATIC1.net" 


.END
