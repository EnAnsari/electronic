** Profile: "SCHEMATIC1-RUN2"  [ C:\Users\WOLF2022\Desktop\UNI\3_semiterm\MadarElectric\Az\word\13\psPise\commonemi-schematic1-run2.sim ] 

** Creating circuit file "commonemi-schematic1-run2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\commonemi-SCHEMATIC1.net" 


.END
