** Profile: "SCHEMATIC1-RUN02"  [ C:\Users\WOLF2022\Desktop\UNI\3_semiterm\MadarElectric\Az\word\13\psPise\commonemi-SCHEMATIC1-RUN02.sim ] 

** Creating circuit file "commonemi-SCHEMATIC1-RUN02.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 1u 
.STEP LIN PARAM RsV 500 2.5k 500 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\commonemi-SCHEMATIC1.net" 


.END
