** Profile: "SCHEMATIC1-RL"  [ C:\Users\WOLF2022\Desktop\UNI\3_semiterm\MadarElectric\Az\word\7-1\RL\rl-schematic1-rl.sim ] 

** Creating circuit file "rl-schematic1-rl.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 1n 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rl-SCHEMATIC1.net" 


.END
