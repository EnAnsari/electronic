** Profile: "SCHEMATIC1-Limit"  [ C:\Users\WOLF2022\Desktop\UNI\3_semiterm\MadarElectric\Az\word\11\Pr0\limiters-schematic1-limit.sim ] 

** Creating circuit file "limiters-schematic1-limit.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\limiters-SCHEMATIC1.net" 


.END
