** Profile: "SCHEMATIC1-RC"  [ C:\Users\WOLF2022\Desktop\UNI\3_semiterm\MadarElectric\Az\word\8\RC\rc-SCHEMATIC1-RC.sim ] 

** Creating circuit file "rc-SCHEMATIC1-RC.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ms 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rc-SCHEMATIC1.net" 


.END
